module orgate
(
    input a,
    input b,
    output x
);

assign x = a | b;

endmodule