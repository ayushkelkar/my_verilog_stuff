module notgate
(
    input a,
    output x
);

assign x = ~a;
endmodule